// ========================================
//  Opcode Table in SPC700 CPU Controller
// ========================================

// Copyright(C) 2024 ep2k All Rights Reserved.

module s_op_table
    import s_cpu_pkg::*;
(
    input logic [7:0] op,

    output addressing_type addressing,
    output instruction_type instruction,
    output reg_src_type reg1_src,
    output reg_src_type reg2_src
);

    addressing_type a;
    instruction_type i;
    reg_src_type r1, r2;

    assign addressing = a;
    assign instruction = i;
    assign reg1_src = r1;
    assign reg2_src = r2;

    always_comb begin
        unique case (op)
            8'h00: {a, i, r1, r2} = {SA_NOP, SI_NOP, SC_R_A, SC_R_A};
            8'h01: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'h02: {a, i, r1, r2} = {SA_SC1_DP, SI_SET1, SC_R_A, SC_R_A};
            8'h03: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBS, SC_R_A, SC_R_A};
            8'h04: {a, i, r1, r2} = {SA_REG_DP, SI_OR, SC_R_A, SC_R_A};
            8'h05: {a, i, r1, r2} = {SA_REG_ABS, SI_OR, SC_R_A, SC_R_A};
            8'h06: {a, i, r1, r2} = {SA_REG_DR, SI_OR, SC_R_A, SC_R_X};
            8'h07: {a, i, r1, r2} = {SA_REG_INDPR, SI_OR, SC_R_A, SC_R_X};
            8'h08: {a, i, r1, r2} = {SA_REG_IMM, SI_OR, SC_R_A, SC_R_A};
            8'h09: {a, i, r1, r2} = {SA_DP_DP, SI_OR, SC_R_A, SC_R_A};
            8'h0A: {a, i, r1, r2} = {SA_CALC1_C_ABS, SI_OR1, SC_R_A, SC_R_A};
            8'h0B: {a, i, r1, r2} = {SA_DP, SI_ASL, SC_R_A, SC_R_A};
            8'h0C: {a, i, r1, r2} = {SA_ABS, SI_ASL, SC_R_A, SC_R_A};
            8'h0D: {a, i, r1, r2} = {SA_PUSH_PSW, SI_PUSH, SC_R_A, SC_R_SP};
            8'h0E: {a, i, r1, r2} = {SA_TSC_ABS, SI_TSET, SC_R_A, SC_R_A};
            8'h0F: {a, i, r1, r2} = {SA_BRK, SI_BRK, SC_R_A, SC_R_A};
            8'h10: {a, i, r1, r2} = {SA_BRA, SI_BPL, SC_R_A, SC_R_A};
            8'h11: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'h12: {a, i, r1, r2} = {SA_SC1_DP, SI_CLR1, SC_R_A, SC_R_A};
            8'h13: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBC, SC_R_A, SC_R_A};
            8'h14: {a, i, r1, r2} = {SA_REG_DPR, SI_OR, SC_R_A, SC_R_X};
            8'h15: {a, i, r1, r2} = {SA_REG_ABSR, SI_OR, SC_R_A, SC_R_X};
            8'h16: {a, i, r1, r2} = {SA_REG_ABSR, SI_OR, SC_R_A, SC_R_Y};
            8'h17: {a, i, r1, r2} = {SA_REG_INDP_R, SI_OR, SC_R_A, SC_R_Y};
            8'h18: {a, i, r1, r2} = {SA_DP_IMM, SI_OR, SC_R_A, SC_R_A};
            8'h19: {a, i, r1, r2} = {SA_DR_DR, SI_OR, SC_R_Y, SC_R_X};
            8'h1A: {a, i, r1, r2} = {SA_DP16, SI_DEC, SC_R_A, SC_R_A};
            8'h1B: {a, i, r1, r2} = {SA_DPR, SI_ASL, SC_R_A, SC_R_X};
            8'h1C: {a, i, r1, r2} = {SA_REG, SI_ASL, SC_R_A, SC_R_A};
            8'h1D: {a, i, r1, r2} = {SA_REG, SI_DEC, SC_R_X, SC_R_A};
            8'h1E: {a, i, r1, r2} = {SA_REG_ABS, SI_CMP, SC_R_X, SC_R_A};
            8'h1F: {a, i, r1, r2} = {SA_JMP_ABSR, SI_JMP, SC_R_A, SC_R_X};
            8'h20: {a, i, r1, r2} = {SA_PSW_CHANGE, SI_CLRP, SC_R_A, SC_R_A};
            8'h21: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'h22: {a, i, r1, r2} = {SA_SC1_DP, SI_SET1, SC_R_A, SC_R_A};
            8'h23: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBS, SC_R_A, SC_R_A};
            8'h24: {a, i, r1, r2} = {SA_REG_DP, SI_AND, SC_R_A, SC_R_A};
            8'h25: {a, i, r1, r2} = {SA_REG_ABS, SI_AND, SC_R_A, SC_R_A};
            8'h26: {a, i, r1, r2} = {SA_REG_DR, SI_AND, SC_R_A, SC_R_X};
            8'h27: {a, i, r1, r2} = {SA_REG_INDPR, SI_AND, SC_R_A, SC_R_X};
            8'h28: {a, i, r1, r2} = {SA_REG_IMM, SI_AND, SC_R_A, SC_R_A};
            8'h29: {a, i, r1, r2} = {SA_DP_DP, SI_AND, SC_R_A, SC_R_A};
            8'h2A: {a, i, r1, r2} = {SA_CALC1_C_ABS, SI_OR1_N, SC_R_A, SC_R_A};
            8'h2B: {a, i, r1, r2} = {SA_DP, SI_ROL, SC_R_A, SC_R_A};
            8'h2C: {a, i, r1, r2} = {SA_ABS, SI_ROL, SC_R_A, SC_R_A};
            8'h2D: {a, i, r1, r2} = {SA_PUSH_REG, SI_PUSH, SC_R_A, SC_R_SP};
            8'h2E: {a, i, r1, r2} = {SA_CBNE_DP, SI_CBNE, SC_R_A, SC_R_A};
            8'h2F: {a, i, r1, r2} = {SA_BRA, SI_BRA, SC_R_A, SC_R_A};
            8'h30: {a, i, r1, r2} = {SA_BRA, SI_BMI, SC_R_A, SC_R_A};
            8'h31: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'h32: {a, i, r1, r2} = {SA_SC1_DP, SI_CLR1, SC_R_A, SC_R_A};
            8'h33: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBC, SC_R_A, SC_R_A};
            8'h34: {a, i, r1, r2} = {SA_REG_DPR, SI_AND, SC_R_A, SC_R_X};
            8'h35: {a, i, r1, r2} = {SA_REG_ABSR, SI_AND, SC_R_A, SC_R_X};
            8'h36: {a, i, r1, r2} = {SA_REG_ABSR, SI_AND, SC_R_A, SC_R_Y};
            8'h37: {a, i, r1, r2} = {SA_REG_INDP_R, SI_AND, SC_R_A, SC_R_Y};
            8'h38: {a, i, r1, r2} = {SA_DP_IMM, SI_AND, SC_R_A, SC_R_A};
            8'h39: {a, i, r1, r2} = {SA_DR_DR, SI_AND, SC_R_Y, SC_R_X};
            8'h3A: {a, i, r1, r2} = {SA_DP16, SI_INC, SC_R_A, SC_R_A};
            8'h3B: {a, i, r1, r2} = {SA_DPR, SI_ROL, SC_R_A, SC_R_X};
            8'h3C: {a, i, r1, r2} = {SA_REG, SI_ROL, SC_R_A, SC_R_A};
            8'h3D: {a, i, r1, r2} = {SA_REG, SI_INC, SC_R_X, SC_R_A};
            8'h3E: {a, i, r1, r2} = {SA_REG_DP, SI_CMP, SC_R_X, SC_R_A};
            8'h3F: {a, i, r1, r2} = {SA_CALL_IMM, SI_CALL, SC_R_A, SC_R_SP};
            8'h40: {a, i, r1, r2} = {SA_PSW_CHANGE, SI_SETP, SC_R_A, SC_R_A};
            8'h41: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'h42: {a, i, r1, r2} = {SA_SC1_DP, SI_SET1, SC_R_A, SC_R_A};
            8'h43: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBS, SC_R_A, SC_R_A};
            8'h44: {a, i, r1, r2} = {SA_REG_DP, SI_EOR, SC_R_A, SC_R_A};
            8'h45: {a, i, r1, r2} = {SA_REG_ABS, SI_EOR, SC_R_A, SC_R_A};
            8'h46: {a, i, r1, r2} = {SA_REG_DR, SI_EOR, SC_R_A, SC_R_X};
            8'h47: {a, i, r1, r2} = {SA_REG_INDPR, SI_EOR, SC_R_A, SC_R_X};
            8'h48: {a, i, r1, r2} = {SA_REG_IMM, SI_EOR, SC_R_A, SC_R_A};
            8'h49: {a, i, r1, r2} = {SA_DP_DP, SI_EOR, SC_R_A, SC_R_A};
            8'h4A: {a, i, r1, r2} = {SA_CALC1_C_ABS, SI_AND1, SC_R_A, SC_R_A};
            8'h4B: {a, i, r1, r2} = {SA_DP, SI_LSR, SC_R_A, SC_R_A};
            8'h4C: {a, i, r1, r2} = {SA_ABS, SI_LSR, SC_R_A, SC_R_A};
            8'h4D: {a, i, r1, r2} = {SA_PUSH_REG, SI_PUSH, SC_R_X, SC_R_SP};
            8'h4E: {a, i, r1, r2} = {SA_TSC_ABS, SI_TCLR, SC_R_A, SC_R_A};
            8'h4F: {a, i, r1, r2} = {SA_CALL_UP, SI_PCALL, SC_R_A, SC_R_SP};
            8'h50: {a, i, r1, r2} = {SA_BRA, SI_BVC, SC_R_A, SC_R_A};
            8'h51: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'h52: {a, i, r1, r2} = {SA_SC1_DP, SI_CLR1, SC_R_A, SC_R_A};
            8'h53: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBC, SC_R_A, SC_R_A};
            8'h54: {a, i, r1, r2} = {SA_REG_DPR, SI_EOR, SC_R_A, SC_R_X};
            8'h55: {a, i, r1, r2} = {SA_REG_ABSR, SI_EOR, SC_R_A, SC_R_X};
            8'h56: {a, i, r1, r2} = {SA_REG_ABSR, SI_EOR, SC_R_A, SC_R_Y};
            8'h57: {a, i, r1, r2} = {SA_REG_INDP_R, SI_EOR, SC_R_A, SC_R_Y};
            8'h58: {a, i, r1, r2} = {SA_DP_IMM, SI_EOR, SC_R_A, SC_R_A};
            8'h59: {a, i, r1, r2} = {SA_DR_DR, SI_EOR, SC_R_Y, SC_R_X};
            8'h5A: {a, i, r1, r2} = {SA_YA_DP16, SI_CMP, SC_R_A, SC_R_Y};
            8'h5B: {a, i, r1, r2} = {SA_DPR, SI_LSR, SC_R_A, SC_R_X};
            8'h5C: {a, i, r1, r2} = {SA_REG, SI_LSR, SC_R_A, SC_R_A};
            8'h5D: {a, i, r1, r2} = {SA_REG_REG, SI_MOV, SC_R_X, SC_R_A};
            8'h5E: {a, i, r1, r2} = {SA_REG_ABS, SI_CMP, SC_R_Y, SC_R_A};
            8'h5F: {a, i, r1, r2} = {SA_JMP_IMM, SI_JMP, SC_R_A, SC_R_A};
            8'h60: {a, i, r1, r2} = {SA_PSW_CHANGE, SI_CLRC, SC_R_A, SC_R_A};
            8'h61: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'h62: {a, i, r1, r2} = {SA_SC1_DP, SI_SET1, SC_R_A, SC_R_A};
            8'h63: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBS, SC_R_A, SC_R_A};
            8'h64: {a, i, r1, r2} = {SA_REG_DP, SI_CMP, SC_R_A, SC_R_A};
            8'h65: {a, i, r1, r2} = {SA_REG_ABS, SI_CMP, SC_R_A, SC_R_A};
            8'h66: {a, i, r1, r2} = {SA_REG_DR, SI_CMP, SC_R_A, SC_R_X};
            8'h67: {a, i, r1, r2} = {SA_REG_INDPR, SI_CMP, SC_R_A, SC_R_X};
            8'h68: {a, i, r1, r2} = {SA_REG_IMM, SI_CMP, SC_R_A, SC_R_A};
            8'h69: {a, i, r1, r2} = {SA_DP_DP, SI_CMP, SC_R_A, SC_R_A};
            8'h6A: {a, i, r1, r2} = {SA_CALC1_C_ABS, SI_AND1_N, SC_R_A, SC_R_A};
            8'h6B: {a, i, r1, r2} = {SA_DP, SI_ROR, SC_R_A, SC_R_A};
            8'h6C: {a, i, r1, r2} = {SA_ABS, SI_ROR, SC_R_A, SC_R_A};
            8'h6D: {a, i, r1, r2} = {SA_PUSH_REG, SI_PUSH, SC_R_Y, SC_R_SP};
            8'h6E: {a, i, r1, r2} = {SA_DBNZ_DP, SI_DBNZ, SC_R_A, SC_R_A};
            8'h6F: {a, i, r1, r2} = {SA_RET, SI_RET, SC_R_A, SC_R_SP};
            8'h70: {a, i, r1, r2} = {SA_BRA, SI_BVS, SC_R_A, SC_R_A};
            8'h71: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'h72: {a, i, r1, r2} = {SA_SC1_DP, SI_CLR1, SC_R_A, SC_R_A};
            8'h73: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBC, SC_R_A, SC_R_A};
            8'h74: {a, i, r1, r2} = {SA_REG_DPR, SI_CMP, SC_R_A, SC_R_X};
            8'h75: {a, i, r1, r2} = {SA_REG_ABSR, SI_CMP, SC_R_A, SC_R_X};
            8'h76: {a, i, r1, r2} = {SA_REG_ABSR, SI_CMP, SC_R_A, SC_R_Y};
            8'h77: {a, i, r1, r2} = {SA_REG_INDP_R, SI_CMP, SC_R_A, SC_R_Y};
            8'h78: {a, i, r1, r2} = {SA_DP_IMM, SI_CMP, SC_R_A, SC_R_A};
            8'h79: {a, i, r1, r2} = {SA_DR_DR, SI_CMP, SC_R_Y, SC_R_X};
            8'h7A: {a, i, r1, r2} = {SA_YA_DP16, SI_ADD, SC_R_A, SC_R_Y};
            8'h7B: {a, i, r1, r2} = {SA_DPR, SI_ROR, SC_R_A, SC_R_X};
            8'h7C: {a, i, r1, r2} = {SA_REG, SI_ROR, SC_R_A, SC_R_A};
            8'h7D: {a, i, r1, r2} = {SA_REG_REG, SI_MOV, SC_R_A, SC_R_X};
            8'h7E: {a, i, r1, r2} = {SA_REG_DP, SI_CMP, SC_R_Y, SC_R_A};
            8'h7F: {a, i, r1, r2} = {SA_RETI, SI_RETI, SC_R_A, SC_R_SP};
            8'h80: {a, i, r1, r2} = {SA_PSW_CHANGE, SI_SETC, SC_R_A, SC_R_A};
            8'h81: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'h82: {a, i, r1, r2} = {SA_SC1_DP, SI_SET1, SC_R_A, SC_R_A};
            8'h83: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBS, SC_R_A, SC_R_A};
            8'h84: {a, i, r1, r2} = {SA_REG_DP, SI_ADC, SC_R_A, SC_R_A};
            8'h85: {a, i, r1, r2} = {SA_REG_ABS, SI_ADC, SC_R_A, SC_R_A};
            8'h86: {a, i, r1, r2} = {SA_REG_DR, SI_ADC, SC_R_A, SC_R_X};
            8'h87: {a, i, r1, r2} = {SA_REG_INDPR, SI_ADC, SC_R_A, SC_R_X};
            8'h88: {a, i, r1, r2} = {SA_REG_IMM, SI_ADC, SC_R_A, SC_R_A};
            8'h89: {a, i, r1, r2} = {SA_DP_DP, SI_ADC, SC_R_A, SC_R_A};
            8'h8A: {a, i, r1, r2} = {SA_CALC1_C_ABS, SI_EOR1, SC_R_A, SC_R_A};
            8'h8B: {a, i, r1, r2} = {SA_DP, SI_DEC, SC_R_A, SC_R_A};
            8'h8C: {a, i, r1, r2} = {SA_ABS, SI_DEC, SC_R_A, SC_R_A};
            8'h8D: {a, i, r1, r2} = {SA_REG_IMM, SI_MOV, SC_R_Y, SC_R_A};
            8'h8E: {a, i, r1, r2} = {SA_POP_PSW, SI_POP, SC_R_A, SC_R_SP};
            8'h8F: {a, i, r1, r2} = {SA_DP_IMM, SI_MOV, SC_R_A, SC_R_A};
            8'h90: {a, i, r1, r2} = {SA_BRA, SI_BCC, SC_R_A, SC_R_A};
            8'h91: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'h92: {a, i, r1, r2} = {SA_SC1_DP, SI_CLR1, SC_R_A, SC_R_A};
            8'h93: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBC, SC_R_A, SC_R_A};
            8'h94: {a, i, r1, r2} = {SA_REG_DPR, SI_ADC, SC_R_A, SC_R_X};
            8'h95: {a, i, r1, r2} = {SA_REG_ABSR, SI_ADC, SC_R_A, SC_R_X};
            8'h96: {a, i, r1, r2} = {SA_REG_ABSR, SI_ADC, SC_R_A, SC_R_Y};
            8'h97: {a, i, r1, r2} = {SA_REG_INDP_R, SI_ADC, SC_R_A, SC_R_Y};
            8'h98: {a, i, r1, r2} = {SA_DP_IMM, SI_ADC, SC_R_A, SC_R_A};
            8'h99: {a, i, r1, r2} = {SA_DR_DR, SI_ADC, SC_R_Y, SC_R_X};
            8'h9A: {a, i, r1, r2} = {SA_YA_DP16, SI_SUB, SC_R_A, SC_R_Y};
            8'h9B: {a, i, r1, r2} = {SA_DPR, SI_DEC, SC_R_A, SC_R_X};
            8'h9C: {a, i, r1, r2} = {SA_REG, SI_DEC, SC_R_A, SC_R_A};
            8'h9D: {a, i, r1, r2} = {SA_REG_REG, SI_MOV, SC_R_X, SC_R_SP};
            8'h9E: {a, i, r1, r2} = {SA_DIV_YA_X, SI_DIV, SC_R_Y, SC_R_X};
            8'h9F: {a, i, r1, r2} = {SA_XCN_REG, SI_XCN, SC_R_A, SC_R_A};
            8'hA0: {a, i, r1, r2} = {SA_PSW_CHANGE, SI_EI, SC_R_A, SC_R_A};
            8'hA1: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'hA2: {a, i, r1, r2} = {SA_SC1_DP, SI_SET1, SC_R_A, SC_R_A};
            8'hA3: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBS, SC_R_A, SC_R_A};
            8'hA4: {a, i, r1, r2} = {SA_REG_DP, SI_SBC, SC_R_A, SC_R_A};
            8'hA5: {a, i, r1, r2} = {SA_REG_ABS, SI_SBC, SC_R_A, SC_R_A};
            8'hA6: {a, i, r1, r2} = {SA_REG_DR, SI_SBC, SC_R_A, SC_R_X};
            8'hA7: {a, i, r1, r2} = {SA_REG_INDPR, SI_SBC, SC_R_A, SC_R_X};
            8'hA8: {a, i, r1, r2} = {SA_REG_IMM, SI_SBC, SC_R_A, SC_R_A};
            8'hA9: {a, i, r1, r2} = {SA_DP_DP, SI_SBC, SC_R_A, SC_R_A};
            8'hAA: {a, i, r1, r2} = {SA_CALC1_C_ABS, SI_MOV1, SC_R_A, SC_R_A};
            8'hAB: {a, i, r1, r2} = {SA_DP, SI_INC, SC_R_A, SC_R_A};
            8'hAC: {a, i, r1, r2} = {SA_ABS, SI_INC, SC_R_A, SC_R_A};
            8'hAD: {a, i, r1, r2} = {SA_REG_IMM, SI_CMP, SC_R_Y, SC_R_A};
            8'hAE: {a, i, r1, r2} = {SA_POP_REG, SI_POP, SC_R_A, SC_R_SP};
            8'hAF: {a, i, r1, r2} = {SA_DRINC_REG, SI_MOV, SC_R_A, SC_R_X};
            8'hB0: {a, i, r1, r2} = {SA_BRA, SI_BCS, SC_R_A, SC_R_A};
            8'hB1: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'hB2: {a, i, r1, r2} = {SA_SC1_DP, SI_CLR1, SC_R_A, SC_R_A};
            8'hB3: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBC, SC_R_A, SC_R_A};
            8'hB4: {a, i, r1, r2} = {SA_REG_DPR, SI_SBC, SC_R_A, SC_R_X};
            8'hB5: {a, i, r1, r2} = {SA_REG_ABSR, SI_SBC, SC_R_A, SC_R_X};
            8'hB6: {a, i, r1, r2} = {SA_REG_ABSR, SI_SBC, SC_R_A, SC_R_Y};
            8'hB7: {a, i, r1, r2} = {SA_REG_INDP_R, SI_SBC, SC_R_A, SC_R_Y};
            8'hB8: {a, i, r1, r2} = {SA_DP_IMM, SI_SBC, SC_R_A, SC_R_A};
            8'hB9: {a, i, r1, r2} = {SA_DR_DR, SI_SBC, SC_R_Y, SC_R_X};
            8'hBA: {a, i, r1, r2} = {SA_YA_DP16, SI_MOV, SC_R_A, SC_R_Y};
            8'hBB: {a, i, r1, r2} = {SA_DPR, SI_INC, SC_R_A, SC_R_X};
            8'hBC: {a, i, r1, r2} = {SA_REG, SI_INC, SC_R_A, SC_R_A};
            8'hBD: {a, i, r1, r2} = {SA_REG_REG, SI_MOV_NF, SC_R_SP, SC_R_X};
            8'hBE: {a, i, r1, r2} = {SA_DAAS, SI_DAS, SC_R_A, SC_R_A};
            8'hBF: {a, i, r1, r2} = {SA_REG_DRINC, SI_MOV, SC_R_A, SC_R_X};
            8'hC0: {a, i, r1, r2} = {SA_PSW_CHANGE, SI_DI, SC_R_A, SC_R_A};
            8'hC1: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'hC2: {a, i, r1, r2} = {SA_SC1_DP, SI_SET1, SC_R_A, SC_R_A};
            8'hC3: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBS, SC_R_A, SC_R_A};
            8'hC4: {a, i, r1, r2} = {SA_DP_REG, SI_MOV, SC_R_A, SC_R_A};
            8'hC5: {a, i, r1, r2} = {SA_ABS_REG, SI_MOV, SC_R_A, SC_R_A};
            8'hC6: {a, i, r1, r2} = {SA_DR_REG, SI_MOV, SC_R_A, SC_R_X};
            8'hC7: {a, i, r1, r2} = {SA_INDPR_REG, SI_MOV, SC_R_A, SC_R_X};
            8'hC8: {a, i, r1, r2} = {SA_REG_IMM, SI_CMP, SC_R_X, SC_R_A};
            8'hC9: {a, i, r1, r2} = {SA_ABS_REG, SI_MOV, SC_R_X, SC_R_A};
            8'hCA: {a, i, r1, r2} = {SA_CALC1_ABS_C, SI_MOV1, SC_R_A, SC_R_A};
            8'hCB: {a, i, r1, r2} = {SA_DP_REG, SI_MOV, SC_R_Y, SC_R_A};
            8'hCC: {a, i, r1, r2} = {SA_ABS_REG, SI_MOV, SC_R_Y, SC_R_A};
            8'hCD: {a, i, r1, r2} = {SA_REG_IMM, SI_MOV, SC_R_X, SC_R_A};
            8'hCE: {a, i, r1, r2} = {SA_POP_REG, SI_POP, SC_R_X, SC_R_SP};
            8'hCF: {a, i, r1, r2} = {SA_MUL_YA, SI_MUL, SC_R_A, SC_R_A};
            8'hD0: {a, i, r1, r2} = {SA_BRA, SI_BNE, SC_R_A, SC_R_A};
            8'hD1: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'hD2: {a, i, r1, r2} = {SA_SC1_DP, SI_CLR1, SC_R_A, SC_R_A};
            8'hD3: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBC, SC_R_A, SC_R_A};
            8'hD4: {a, i, r1, r2} = {SA_DPR_REG, SI_MOV, SC_R_A, SC_R_X};
            8'hD5: {a, i, r1, r2} = {SA_ABSR_REG, SI_MOV, SC_R_A, SC_R_X};
            8'hD6: {a, i, r1, r2} = {SA_ABSR_REG, SI_MOV, SC_R_A, SC_R_Y};
            8'hD7: {a, i, r1, r2} = {SA_INDP_R_REG, SI_MOV, SC_R_A, SC_R_Y};
            8'hD8: {a, i, r1, r2} = {SA_DP_REG, SI_MOV, SC_R_X, SC_R_A};
            8'hD9: {a, i, r1, r2} = {SA_DPR_REG, SI_MOV, SC_R_X, SC_R_Y};
            8'hDA: {a, i, r1, r2} = {SA_DP16_YA, SI_MOV, SC_R_A, SC_R_Y};
            8'hDB: {a, i, r1, r2} = {SA_DPR_REG, SI_MOV, SC_R_Y, SC_R_X};
            8'hDC: {a, i, r1, r2} = {SA_REG, SI_DEC, SC_R_Y, SC_R_A};
            8'hDD: {a, i, r1, r2} = {SA_REG_REG, SI_MOV, SC_R_A, SC_R_Y};
            8'hDE: {a, i, r1, r2} = {SA_CBNE_DPR, SI_CBNE, SC_R_A, SC_R_X};
            8'hDF: {a, i, r1, r2} = {SA_DAAS, SI_DAA, SC_R_A, SC_R_A};
            8'hE0: {a, i, r1, r2} = {SA_PSW_CHANGE, SI_CLRV, SC_R_A, SC_R_A};
            8'hE1: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'hE2: {a, i, r1, r2} = {SA_SC1_DP, SI_SET1, SC_R_A, SC_R_A};
            8'hE3: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBS, SC_R_A, SC_R_A};
            8'hE4: {a, i, r1, r2} = {SA_REG_DP, SI_MOV, SC_R_A, SC_R_A};
            8'hE5: {a, i, r1, r2} = {SA_REG_ABS, SI_MOV, SC_R_A, SC_R_A};
            8'hE6: {a, i, r1, r2} = {SA_REG_DR, SI_MOV, SC_R_A, SC_R_X};
            8'hE7: {a, i, r1, r2} = {SA_REG_INDPR, SI_MOV, SC_R_A, SC_R_X};
            8'hE8: {a, i, r1, r2} = {SA_REG_IMM, SI_MOV, SC_R_A, SC_R_A};
            8'hE9: {a, i, r1, r2} = {SA_REG_ABS, SI_MOV, SC_R_X, SC_R_A};
            8'hEA: {a, i, r1, r2} = {SA_CALC1_ABS_C, SI_NOT1, SC_R_A, SC_R_A};
            8'hEB: {a, i, r1, r2} = {SA_REG_DP, SI_MOV, SC_R_Y, SC_R_A};
            8'hEC: {a, i, r1, r2} = {SA_REG_ABS, SI_MOV, SC_R_Y, SC_R_A};
            8'hED: {a, i, r1, r2} = {SA_PSW_CHANGE, SI_NOTC, SC_R_A, SC_R_A};
            8'hEE: {a, i, r1, r2} = {SA_POP_REG, SI_POP, SC_R_Y, SC_R_SP};
            8'hEF: {a, i, r1, r2} = {SA_NOP, SI_SLEEP, SC_R_A, SC_R_A};
            8'hF0: {a, i, r1, r2} = {SA_BRA, SI_BEQ, SC_R_A, SC_R_A};
            8'hF1: {a, i, r1, r2} = {SA_CALL_N, SI_TCALL, SC_R_A, SC_R_SP};
            8'hF2: {a, i, r1, r2} = {SA_SC1_DP, SI_CLR1, SC_R_A, SC_R_A};
            8'hF3: {a, i, r1, r2} = {SA_BBSC_DP, SI_BBC, SC_R_A, SC_R_A};
            8'hF4: {a, i, r1, r2} = {SA_REG_DPR, SI_MOV, SC_R_A, SC_R_X};
            8'hF5: {a, i, r1, r2} = {SA_REG_ABSR, SI_MOV, SC_R_A, SC_R_X};
            8'hF6: {a, i, r1, r2} = {SA_REG_ABSR, SI_MOV, SC_R_A, SC_R_Y};
            8'hF7: {a, i, r1, r2} = {SA_REG_INDP_R, SI_MOV, SC_R_A, SC_R_Y};
            8'hF8: {a, i, r1, r2} = {SA_REG_DP, SI_MOV, SC_R_X, SC_R_A};
            8'hF9: {a, i, r1, r2} = {SA_REG_DPR, SI_MOV, SC_R_X, SC_R_Y};
            8'hFA: {a, i, r1, r2} = {SA_DP_DP, SI_MOV, SC_R_A, SC_R_A};
            8'hFB: {a, i, r1, r2} = {SA_REG_DPR, SI_MOV, SC_R_Y, SC_R_X};
            8'hFC: {a, i, r1, r2} = {SA_REG, SI_INC, SC_R_Y, SC_R_A};
            8'hFD: {a, i, r1, r2} = {SA_REG_REG, SI_MOV, SC_R_Y, SC_R_A};
            8'hFE: {a, i, r1, r2} = {SA_DBNZ_REG, SI_DBNZ, SC_R_A, SC_R_Y};
            8'hFF: {a, i, r1, r2} = {SA_NOP, SI_STOP, SC_R_A, SC_R_A};
        endcase
    end
    
endmodule
