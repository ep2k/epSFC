// ========================================
//  Opecode Table in 65816 CPU Controller
// ========================================

// Copyright(C) 2024 ep2k All Rights Reserved.

module opcode_table
    import cpu_pkg::*;
(
    input logic [7:0] op,
    input logic m8,

    output addressing_type addressing,
    output instruction_type instruction,
    output logic [2:0] init_op_counter
);

    always_comb begin
        unique case (op)
            8'h00: {addressing, instruction} = {A_SOFT_INT, I_BRK};
            8'h01: {addressing, instruction} = {A_INDPX, I_ORA};
            8'h02: {addressing, instruction} = {A_SOFT_INT, I_COP};
            8'h03: {addressing, instruction} = {A_SPR, I_ORA};
            8'h04: {addressing, instruction} = {A_DP, I_TSB};
            8'h05: {addressing, instruction} = {A_DP, I_ORA};
            8'h06: {addressing, instruction} = {A_DP, I_ASL};
            8'h07: {addressing, instruction} = {A_INDPL, I_ORA};
            8'h08: {addressing, instruction} = {A_PUSH_P, I_PHA};
            8'h09: {addressing, instruction} = {A_IMM, I_ORA};
            8'h0A: {addressing, instruction} = {A_IMP, I_ASL_A};
            8'h0B: {addressing, instruction} = {A_PUSH_DP, I_PHA};
            8'h0C: {addressing, instruction} = {A_ABS, I_TSB};
            8'h0D: {addressing, instruction} = {A_ABS, I_ORA};
            8'h0E: {addressing, instruction} = {A_ABS, I_ASL};
            8'h0F: {addressing, instruction} = {A_ABSL, I_ORA};
            8'h10: {addressing, instruction} = {A_IMP, I_BPL};
            8'h11: {addressing, instruction} = {A_INDPY, I_ORA};
            8'h12: {addressing, instruction} = {A_INDP, I_ORA};
            8'h13: {addressing, instruction} = {A_INSPRY, I_ORA};
            8'h14: {addressing, instruction} = {A_DP, I_TRB};
            8'h15: {addressing, instruction} = {A_DPX, I_ORA};
            8'h16: {addressing, instruction} = {A_DPX, I_ASL};
            8'h17: {addressing, instruction} = {A_INDPLY, I_ORA};
            8'h18: {addressing, instruction} = {A_IMP, I_CLC};
            8'h19: {addressing, instruction} = {A_ABSY, I_ORA};
            8'h1A: {addressing, instruction} = {A_IMP, I_INC_A};
            8'h1B: {addressing, instruction} = {A_IMP, I_TCS};
            8'h1C: {addressing, instruction} = {A_ABS, I_TRB};
            8'h1D: {addressing, instruction} = {A_ABSX, I_ORA};
            8'h1E: {addressing, instruction} = {A_ABSX, I_ASL};
            8'h1F: {addressing, instruction} = {A_ABSLX, I_ORA};
            8'h20: {addressing, instruction} = {A_SUB_IMM, I_JSR};
            8'h21: {addressing, instruction} = {A_INDPX, I_AND};
            8'h22: {addressing, instruction} = {A_SUB_IMML, I_JSR};
            8'h23: {addressing, instruction} = {A_SPR, I_AND};
            8'h24: {addressing, instruction} = {A_DP, I_BIT};
            8'h25: {addressing, instruction} = {A_DP, I_AND};
            8'h26: {addressing, instruction} = {A_DP, I_ROL};
            8'h27: {addressing, instruction} = {A_INDPL, I_AND};
            8'h28: {addressing, instruction} = {A_PULL_P, I_PLA};
            8'h29: {addressing, instruction} = {A_IMM, I_AND};
            8'h2A: {addressing, instruction} = {A_IMP, I_ROL_A};
            8'h2B: {addressing, instruction} = {A_PULL_DP, I_PLA};
            8'h2C: {addressing, instruction} = {A_ABS, I_BIT};
            8'h2D: {addressing, instruction} = {A_ABS, I_AND};
            8'h2E: {addressing, instruction} = {A_ABS, I_ROL};
            8'h2F: {addressing, instruction} = {A_ABSL, I_AND};
            8'h30: {addressing, instruction} = {A_IMP, I_BMI};
            8'h31: {addressing, instruction} = {A_INDPY, I_AND};
            8'h32: {addressing, instruction} = {A_INDP, I_AND};
            8'h33: {addressing, instruction} = {A_INSPRY, I_AND};
            8'h34: {addressing, instruction} = {A_DPX, I_BIT};
            8'h35: {addressing, instruction} = {A_DPX, I_AND};
            8'h36: {addressing, instruction} = {A_DPX, I_ROL};
            8'h37: {addressing, instruction} = {A_INDPLY, I_AND};
            8'h38: {addressing, instruction} = {A_IMP, I_SEC};
            8'h39: {addressing, instruction} = {A_ABSY, I_AND};
            8'h3A: {addressing, instruction} = {A_IMP, I_DEC_A};
            8'h3B: {addressing, instruction} = {A_IMP, I_TSC};
            8'h3C: {addressing, instruction} = {A_ABSX, I_BIT};
            8'h3D: {addressing, instruction} = {A_ABSX, I_AND};
            8'h3E: {addressing, instruction} = {A_ABSX, I_ROL};
            8'h3F: {addressing, instruction} = {A_ABSLX, I_AND};
            8'h40: {addressing, instruction} = {A_RTI, I_RTI};
            8'h41: {addressing, instruction} = {A_INDPX, I_EOR};
            8'h42: {addressing, instruction} = {A_IMP, I_WDM};
            8'h43: {addressing, instruction} = {A_SPR, I_EOR};
            8'h44: {addressing, instruction} = {A_MVP, I_MVP};
            8'h45: {addressing, instruction} = {A_DP, I_EOR};
            8'h46: {addressing, instruction} = {A_DP, I_LSR};
            8'h47: {addressing, instruction} = {A_INDPL, I_EOR};
            8'h48: {addressing, instruction} = {A_PUSH_A, I_PHA};
            8'h49: {addressing, instruction} = {A_IMM, I_EOR};
            8'h4A: {addressing, instruction} = {A_IMP, I_LSR_A};
            8'h4B: {addressing, instruction} = {A_PUSH_PB, I_PHA};
            8'h4C: {addressing, instruction} = {A_IMM_JMP, I_JMP};
            8'h4D: {addressing, instruction} = {A_ABS, I_EOR};
            8'h4E: {addressing, instruction} = {A_ABS, I_LSR};
            8'h4F: {addressing, instruction} = {A_ABSL, I_EOR};
            8'h50: {addressing, instruction} = {A_IMP, I_BVC};
            8'h51: {addressing, instruction} = {A_INDPY, I_EOR};
            8'h52: {addressing, instruction} = {A_INDP, I_EOR};
            8'h53: {addressing, instruction} = {A_INSPRY, I_EOR};
            8'h54: {addressing, instruction} = {A_MVN, I_MVN};
            8'h55: {addressing, instruction} = {A_DPX, I_EOR};
            8'h56: {addressing, instruction} = {A_DPX, I_LSR};
            8'h57: {addressing, instruction} = {A_INDPLY, I_EOR};
            8'h58: {addressing, instruction} = {A_IMP, I_CLI};
            8'h59: {addressing, instruction} = {A_ABSY, I_EOR};
            8'h5A: {addressing, instruction} = {A_PUSH_Y, I_PHA};
            8'h5B: {addressing, instruction} = {A_IMP, I_TCD};
            8'h5C: {addressing, instruction} = {A_IMM_JMP, I_JMPL};
            8'h5D: {addressing, instruction} = {A_ABSX, I_EOR};
            8'h5E: {addressing, instruction} = {A_ABSX, I_LSR};
            8'h5F: {addressing, instruction} = {A_ABSLX, I_EOR};
            8'h60: {addressing, instruction} = {A_RTS, I_RTS};
            8'h61: {addressing, instruction} = {A_INDPX, I_ADC};
            8'h62: {addressing, instruction} = {A_PER, I_PER};
            8'h63: {addressing, instruction} = {A_SPR, I_ADC};
            8'h64: {addressing, instruction} = {A_DP, I_STZ};
            8'h65: {addressing, instruction} = {A_DP, I_ADC};
            8'h66: {addressing, instruction} = {A_DP, I_ROR};
            8'h67: {addressing, instruction} = {A_INDPL, I_ADC};
            8'h68: {addressing, instruction} = {A_PULL_A, I_PLA};
            8'h69: {addressing, instruction} = {A_IMM, I_ADC};
            8'h6A: {addressing, instruction} = {A_IMP, I_ROR_A};
            8'h6B: {addressing, instruction} = {A_RTL, I_RTL};
            8'h6C: {addressing, instruction} = {A_ABS_JMP, I_JMP};
            8'h6D: {addressing, instruction} = {A_ABS, I_ADC};
            8'h6E: {addressing, instruction} = {A_ABS, I_ROR};
            8'h6F: {addressing, instruction} = {A_ABSL, I_ADC};
            8'h70: {addressing, instruction} = {A_IMP, I_BVS};
            8'h71: {addressing, instruction} = {A_INDPY, I_ADC};
            8'h72: {addressing, instruction} = {A_INDP, I_ADC};
            8'h73: {addressing, instruction} = {A_INSPRY, I_ADC};
            8'h74: {addressing, instruction} = {A_DPX, I_STZ};
            8'h75: {addressing, instruction} = {A_DPX, I_ADC};
            8'h76: {addressing, instruction} = {A_DPX, I_ROR};
            8'h77: {addressing, instruction} = {A_INDPLY, I_ADC};
            8'h78: {addressing, instruction} = {A_IMP, I_SEI};
            8'h79: {addressing, instruction} = {A_ABSY, I_ADC};
            8'h7A: {addressing, instruction} = {A_PULL_Y, I_PLA};
            8'h7B: {addressing, instruction} = {A_IMP, I_TDC};
            8'h7C: {addressing, instruction} = {A_ABSX_JMP, I_JMP};
            8'h7D: {addressing, instruction} = {A_ABSX, I_ADC};
            8'h7E: {addressing, instruction} = {A_ABSX, I_ROR};
            8'h7F: {addressing, instruction} = {A_ABSLX, I_ADC};
            8'h80: {addressing, instruction} = {A_IMP, I_BRA};
            8'h81: {addressing, instruction} = {A_INDPX, I_STA};
            8'h82: {addressing, instruction} = {A_IMP, I_BRL};
            8'h83: {addressing, instruction} = {A_SPR, I_STA};
            8'h84: {addressing, instruction} = {A_DP, I_STY};
            8'h85: {addressing, instruction} = {A_DP, I_STA};
            8'h86: {addressing, instruction} = {A_DP, I_STX};
            8'h87: {addressing, instruction} = {A_INDPL, I_STA};
            8'h88: {addressing, instruction} = {A_IMP, I_DEY};
            8'h89: {addressing, instruction} = {A_IMM, I_BIT};
            8'h8A: {addressing, instruction} = {A_IMP, I_TXA};
            8'h8B: {addressing, instruction} = {A_PUSH_DB, I_PHA};
            8'h8C: {addressing, instruction} = {A_ABS, I_STY};
            8'h8D: {addressing, instruction} = {A_ABS, I_STA};
            8'h8E: {addressing, instruction} = {A_ABS, I_STX};
            8'h8F: {addressing, instruction} = {A_ABSL, I_STA};
            8'h90: {addressing, instruction} = {A_IMP, I_BCC};
            8'h91: {addressing, instruction} = {A_INDPY, I_STA};
            8'h92: {addressing, instruction} = {A_INDP, I_STA};
            8'h93: {addressing, instruction} = {A_INSPRY, I_STA};
            8'h94: {addressing, instruction} = {A_DPX, I_STY};
            8'h95: {addressing, instruction} = {A_DPX, I_STA};
            8'h96: {addressing, instruction} = {A_DPY, I_STX};
            8'h97: {addressing, instruction} = {A_INDPLY, I_STA};
            8'h98: {addressing, instruction} = {A_IMP, I_TYA};
            8'h99: {addressing, instruction} = {A_ABSY, I_STA};
            8'h9A: {addressing, instruction} = {A_IMP, I_TXS};
            8'h9B: {addressing, instruction} = {A_IMP, I_TXY};
            8'h9C: {addressing, instruction} = {A_ABS, I_STZ};
            8'h9D: {addressing, instruction} = {A_ABSX, I_STA};
            8'h9E: {addressing, instruction} = {A_ABSX, I_STZ};
            8'h9F: {addressing, instruction} = {A_ABSLX, I_STA};
            8'hA0: {addressing, instruction} = {A_IMM, I_LDY};
            8'hA1: {addressing, instruction} = {A_INDPX, I_LDA};
            8'hA2: {addressing, instruction} = {A_IMM, I_LDX};
            8'hA3: {addressing, instruction} = {A_SPR, I_LDA};
            8'hA4: {addressing, instruction} = {A_DP, I_LDY};
            8'hA5: {addressing, instruction} = {A_DP, I_LDA};
            8'hA6: {addressing, instruction} = {A_DP, I_LDX};
            8'hA7: {addressing, instruction} = {A_INDPL, I_LDA};
            8'hA8: {addressing, instruction} = {A_IMP, I_TAY};
            8'hA9: {addressing, instruction} = {A_IMM, I_LDA};
            8'hAA: {addressing, instruction} = {A_IMP, I_TAX};
            8'hAB: {addressing, instruction} = {A_PULL_DB, I_PLA};
            8'hAC: {addressing, instruction} = {A_ABS, I_LDY};
            8'hAD: {addressing, instruction} = {A_ABS, I_LDA};
            8'hAE: {addressing, instruction} = {A_ABS, I_LDX};
            8'hAF: {addressing, instruction} = {A_ABSL, I_LDA};
            8'hB0: {addressing, instruction} = {A_IMP, I_BCS};
            8'hB1: {addressing, instruction} = {A_INDPY, I_LDA};
            8'hB2: {addressing, instruction} = {A_INDP, I_LDA};
            8'hB3: {addressing, instruction} = {A_INSPRY, I_LDA};
            8'hB4: {addressing, instruction} = {A_DPX, I_LDY};
            8'hB5: {addressing, instruction} = {A_DPX, I_LDA};
            8'hB6: {addressing, instruction} = {A_DPY, I_LDX};
            8'hB7: {addressing, instruction} = {A_INDPLY, I_LDA};
            8'hB8: {addressing, instruction} = {A_IMP, I_CLV};
            8'hB9: {addressing, instruction} = {A_ABSY, I_LDA};
            8'hBA: {addressing, instruction} = {A_IMP, I_TSX};
            8'hBB: {addressing, instruction} = {A_IMP, I_TYX};
            8'hBC: {addressing, instruction} = {A_ABSX, I_LDY};
            8'hBD: {addressing, instruction} = {A_ABSX, I_LDA};
            8'hBE: {addressing, instruction} = {A_ABSY, I_LDX};
            8'hBF: {addressing, instruction} = {A_ABSLX, I_LDA};
            8'hC0: {addressing, instruction} = {A_IMM, I_CPY};
            8'hC1: {addressing, instruction} = {A_INDPX, I_CMP};
            8'hC2: {addressing, instruction} = {A_IMM, I_REP};
            8'hC3: {addressing, instruction} = {A_SPR, I_CMP};
            8'hC4: {addressing, instruction} = {A_DP, I_CPY};
            8'hC5: {addressing, instruction} = {A_DP, I_CMP};
            8'hC6: {addressing, instruction} = {A_DP, I_DEC};
            8'hC7: {addressing, instruction} = {A_INDPL, I_CMP};
            8'hC8: {addressing, instruction} = {A_IMP, I_INY};
            8'hC9: {addressing, instruction} = {A_IMM, I_CMP};
            8'hCA: {addressing, instruction} = {A_IMP, I_DEX};
            8'hCB: {addressing, instruction} = {A_WAIT, I_WAI};
            8'hCC: {addressing, instruction} = {A_ABS, I_CPY};
            8'hCD: {addressing, instruction} = {A_ABS, I_CMP};
            8'hCE: {addressing, instruction} = {A_ABS, I_DEC};
            8'hCF: {addressing, instruction} = {A_ABSL, I_CMP};
            8'hD0: {addressing, instruction} = {A_IMP, I_BNE};
            8'hD1: {addressing, instruction} = {A_INDPY, I_CMP};
            8'hD2: {addressing, instruction} = {A_INDP, I_CMP};
            8'hD3: {addressing, instruction} = {A_INSPRY, I_CMP};
            8'hD4: {addressing, instruction} = {A_PEI, I_PEI};
            8'hD5: {addressing, instruction} = {A_DPX, I_CMP};
            8'hD6: {addressing, instruction} = {A_DPX, I_DEC};
            8'hD7: {addressing, instruction} = {A_INDPLY, I_CMP};
            8'hD8: {addressing, instruction} = {A_IMP, I_CLD};
            8'hD9: {addressing, instruction} = {A_ABSY, I_CMP};
            8'hDA: {addressing, instruction} = {A_PUSH_X, I_PHA};
            8'hDB: {addressing, instruction} = {A_WAIT, I_STP};
            8'hDC: {addressing, instruction} = {A_ABSL_JMP, I_JMPL};
            8'hDD: {addressing, instruction} = {A_ABSX, I_CMP};
            8'hDE: {addressing, instruction} = {A_ABSX, I_DEC};
            8'hDF: {addressing, instruction} = {A_ABSLX, I_CMP};
            8'hE0: {addressing, instruction} = {A_IMM, I_CPX};
            8'hE1: {addressing, instruction} = {A_INDPX, I_SBC};
            8'hE2: {addressing, instruction} = {A_IMM, I_SEP};
            8'hE3: {addressing, instruction} = {A_SPR, I_SBC};
            8'hE4: {addressing, instruction} = {A_DP, I_CPX};
            8'hE5: {addressing, instruction} = {A_DP, I_SBC};
            8'hE6: {addressing, instruction} = {A_DP, I_INC};
            8'hE7: {addressing, instruction} = {A_INDPL, I_SBC};
            8'hE8: {addressing, instruction} = {A_IMP, I_INX};
            8'hE9: {addressing, instruction} = {A_IMM, I_SBC};
            8'hEA: {addressing, instruction} = {A_IMP, I_NOP};
            8'hEB: {addressing, instruction} = {A_IMP, I_XBA};
            8'hEC: {addressing, instruction} = {A_ABS, I_CPX};
            8'hED: {addressing, instruction} = {A_ABS, I_SBC};
            8'hEE: {addressing, instruction} = {A_ABS, I_INC};
            8'hEF: {addressing, instruction} = {A_ABSL, I_SBC};
            8'hF0: {addressing, instruction} = {A_IMP, I_BEQ};
            8'hF1: {addressing, instruction} = {A_INDPY, I_SBC};
            8'hF2: {addressing, instruction} = {A_INDP, I_SBC};
            8'hF3: {addressing, instruction} = {A_INSPRY, I_SBC};
            8'hF4: {addressing, instruction} = {A_PEA, I_PEA};
            8'hF5: {addressing, instruction} = {A_DPX, I_SBC};
            8'hF6: {addressing, instruction} = {A_DPX, I_INC};
            8'hF7: {addressing, instruction} = {A_INDPLY, I_SBC};
            8'hF8: {addressing, instruction} = {A_IMP, I_SED};
            8'hF9: {addressing, instruction} = {A_ABSY, I_SBC};
            8'hFA: {addressing, instruction} = {A_PULL_X, I_PLA};
            8'hFB: {addressing, instruction} = {A_IMP, I_XCE};
            8'hFC: {addressing, instruction} = {A_SUB_ABSX, I_JSR};
            8'hFD: {addressing, instruction} = {A_ABSX, I_SBC};
            8'hFE: {addressing, instruction} = {A_ABSX, I_INC};
            8'hFF: {addressing, instruction} = {A_ABSLX, I_SBC};
        endcase
    end

    always_comb begin
        case (instruction)
            I_LDA: init_op_counter = 3'd1;
            I_LDX: init_op_counter = 3'd1;
            I_LDY: init_op_counter = 3'd1;
            I_STA: init_op_counter = 3'd1;
            I_STX: init_op_counter = 3'd1;
            I_STY: init_op_counter = 3'd1;
            I_STZ: init_op_counter = 3'd1;
            I_ADC: init_op_counter = 3'd1;
            I_SBC: init_op_counter = 3'd1;
            I_AND: init_op_counter = 3'd1;
            I_EOR: init_op_counter = 3'd1;
            I_ORA: init_op_counter = 3'd1;
            I_BIT: init_op_counter = 3'd1;
            I_REP: init_op_counter = 3'd1;
            I_SEP: init_op_counter = 3'd1;
            I_CMP: init_op_counter = 3'd1;
            I_CPX: init_op_counter = 3'd1;
            I_CPY: init_op_counter = 3'd1;
            I_INC_A: init_op_counter = 3'd0;
            I_DEC_A: init_op_counter = 3'd0;
            I_ASL_A: init_op_counter = 3'd0;
            I_LSR_A: init_op_counter = 3'd0;
            I_ROL_A: init_op_counter = 3'd0;
            I_ROR_A: init_op_counter = 3'd0;
            I_INX: init_op_counter = 3'd0;
            I_INY: init_op_counter = 3'd0;
            I_DEX: init_op_counter = 3'd0;
            I_DEY: init_op_counter = 3'd0;
            I_INC: init_op_counter = 3'd4 - m8;
            I_DEC: init_op_counter = 3'd4 - m8;
            I_ASL: init_op_counter = 3'd4 - m8;
            I_LSR: init_op_counter = 3'd4 - m8;
            I_ROL: init_op_counter = 3'd4 - m8;
            I_ROR: init_op_counter = 3'd4 - m8;
            I_TRB: init_op_counter = 3'd4 - m8;
            I_TSB: init_op_counter = 3'd4 - m8;
            I_BCC: init_op_counter = 3'd2;
            I_BCS: init_op_counter = 3'd2;
            I_BEQ: init_op_counter = 3'd2;
            I_BMI: init_op_counter = 3'd2;
            I_BNE: init_op_counter = 3'd2;
            I_BPL: init_op_counter = 3'd2;
            I_BRA: init_op_counter = 3'd2;
            I_BVC: init_op_counter = 3'd2;
            I_BVS: init_op_counter = 3'd2;
            I_BRL: init_op_counter = 3'd2;
            I_JMP: init_op_counter = 3'd2;
            I_JMPL: init_op_counter = 3'd2;
            I_CLC: init_op_counter = 3'd0;
            I_CLD: init_op_counter = 3'd0;
            I_CLI: init_op_counter = 3'd0;
            I_CLV: init_op_counter = 3'd0;
            I_SEC: init_op_counter = 3'd0;
            I_SED: init_op_counter = 3'd0;
            I_SEI: init_op_counter = 3'd0;
            I_TAX: init_op_counter = 3'd0;
            I_TAY: init_op_counter = 3'd0;
            I_TSX: init_op_counter = 3'd0;
            I_TXA: init_op_counter = 3'd0;
            I_TXS: init_op_counter = 3'd0;
            I_TXY: init_op_counter = 3'd0;
            I_TYA: init_op_counter = 3'd0;
            I_TYX: init_op_counter = 3'd0;
            I_TCD: init_op_counter = 3'd0;
            I_TCS: init_op_counter = 3'd0;
            I_TDC: init_op_counter = 3'd0;
            I_TSC: init_op_counter = 3'd0;
            I_PHA: init_op_counter = 3'd0;
            I_PLA: init_op_counter = 3'd1;
            I_RTI: init_op_counter = 3'd1;
            I_RTL: init_op_counter = 3'd1;
            I_RTS: init_op_counter = 3'd2;
            I_XBA: init_op_counter = 3'd1;
            I_XCE: init_op_counter = 3'd0;
            I_BRK: init_op_counter = 3'd1;
            I_COP: init_op_counter = 3'd1;
            default: init_op_counter = 3'd0;
        endcase
    end
    
endmodule
