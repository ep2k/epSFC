// ==============================
//  Brightness Table
// ==============================

// Copyright(C) 2024 ep2k All Rights Reserved.

module brightness_table (
    input logic [4:0] color_raw,
    input logic [3:0] brightness,

    output logic [4:0] color
);

    // color = color_raw * (brightness + 1) / 16
    // brightness = 0 の場合は color = 0
    // [TODO] 乗算器を使うべきか
    always_comb begin
        case ({brightness, color_raw})
            {4'h1, 5'h0}: color = 5'h0;
            {4'h1, 5'h1}: color = 5'h0;
            {4'h1, 5'h2}: color = 5'h0;
            {4'h1, 5'h3}: color = 5'h0;
            {4'h1, 5'h4}: color = 5'h1;
            {4'h1, 5'h5}: color = 5'h1;
            {4'h1, 5'h6}: color = 5'h1;
            {4'h1, 5'h7}: color = 5'h1;
            {4'h1, 5'h8}: color = 5'h1;
            {4'h1, 5'h9}: color = 5'h1;
            {4'h1, 5'hA}: color = 5'h1;
            {4'h1, 5'hB}: color = 5'h1;
            {4'h1, 5'hC}: color = 5'h2;
            {4'h1, 5'hD}: color = 5'h2;
            {4'h1, 5'hE}: color = 5'h2;
            {4'h1, 5'hF}: color = 5'h2;
            {4'h1, 5'h10}: color = 5'h2;
            {4'h1, 5'h11}: color = 5'h2;
            {4'h1, 5'h12}: color = 5'h2;
            {4'h1, 5'h13}: color = 5'h2;
            {4'h1, 5'h14}: color = 5'h3;
            {4'h1, 5'h15}: color = 5'h3;
            {4'h1, 5'h16}: color = 5'h3;
            {4'h1, 5'h17}: color = 5'h3;
            {4'h1, 5'h18}: color = 5'h3;
            {4'h1, 5'h19}: color = 5'h3;
            {4'h1, 5'h1A}: color = 5'h3;
            {4'h1, 5'h1B}: color = 5'h3;
            {4'h1, 5'h1C}: color = 5'h4;
            {4'h1, 5'h1D}: color = 5'h4;
            {4'h1, 5'h1E}: color = 5'h4;
            {4'h1, 5'h1F}: color = 5'h4;
            {4'h2, 5'h0}: color = 5'h0;
            {4'h2, 5'h1}: color = 5'h0;
            {4'h2, 5'h2}: color = 5'h0;
            {4'h2, 5'h3}: color = 5'h1;
            {4'h2, 5'h4}: color = 5'h1;
            {4'h2, 5'h5}: color = 5'h1;
            {4'h2, 5'h6}: color = 5'h1;
            {4'h2, 5'h7}: color = 5'h1;
            {4'h2, 5'h8}: color = 5'h2;
            {4'h2, 5'h9}: color = 5'h2;
            {4'h2, 5'hA}: color = 5'h2;
            {4'h2, 5'hB}: color = 5'h2;
            {4'h2, 5'hC}: color = 5'h2;
            {4'h2, 5'hD}: color = 5'h2;
            {4'h2, 5'hE}: color = 5'h3;
            {4'h2, 5'hF}: color = 5'h3;
            {4'h2, 5'h10}: color = 5'h3;
            {4'h2, 5'h11}: color = 5'h3;
            {4'h2, 5'h12}: color = 5'h3;
            {4'h2, 5'h13}: color = 5'h4;
            {4'h2, 5'h14}: color = 5'h4;
            {4'h2, 5'h15}: color = 5'h4;
            {4'h2, 5'h16}: color = 5'h4;
            {4'h2, 5'h17}: color = 5'h4;
            {4'h2, 5'h18}: color = 5'h5;
            {4'h2, 5'h19}: color = 5'h5;
            {4'h2, 5'h1A}: color = 5'h5;
            {4'h2, 5'h1B}: color = 5'h5;
            {4'h2, 5'h1C}: color = 5'h5;
            {4'h2, 5'h1D}: color = 5'h5;
            {4'h2, 5'h1E}: color = 5'h6;
            {4'h2, 5'h1F}: color = 5'h6;
            {4'h3, 5'h0}: color = 5'h0;
            {4'h3, 5'h1}: color = 5'h0;
            {4'h3, 5'h2}: color = 5'h1;
            {4'h3, 5'h3}: color = 5'h1;
            {4'h3, 5'h4}: color = 5'h1;
            {4'h3, 5'h5}: color = 5'h1;
            {4'h3, 5'h6}: color = 5'h2;
            {4'h3, 5'h7}: color = 5'h2;
            {4'h3, 5'h8}: color = 5'h2;
            {4'h3, 5'h9}: color = 5'h2;
            {4'h3, 5'hA}: color = 5'h3;
            {4'h3, 5'hB}: color = 5'h3;
            {4'h3, 5'hC}: color = 5'h3;
            {4'h3, 5'hD}: color = 5'h3;
            {4'h3, 5'hE}: color = 5'h4;
            {4'h3, 5'hF}: color = 5'h4;
            {4'h3, 5'h10}: color = 5'h4;
            {4'h3, 5'h11}: color = 5'h4;
            {4'h3, 5'h12}: color = 5'h5;
            {4'h3, 5'h13}: color = 5'h5;
            {4'h3, 5'h14}: color = 5'h5;
            {4'h3, 5'h15}: color = 5'h5;
            {4'h3, 5'h16}: color = 5'h6;
            {4'h3, 5'h17}: color = 5'h6;
            {4'h3, 5'h18}: color = 5'h6;
            {4'h3, 5'h19}: color = 5'h6;
            {4'h3, 5'h1A}: color = 5'h7;
            {4'h3, 5'h1B}: color = 5'h7;
            {4'h3, 5'h1C}: color = 5'h7;
            {4'h3, 5'h1D}: color = 5'h7;
            {4'h3, 5'h1E}: color = 5'h8;
            {4'h3, 5'h1F}: color = 5'h8;
            {4'h4, 5'h0}: color = 5'h0;
            {4'h4, 5'h1}: color = 5'h0;
            {4'h4, 5'h2}: color = 5'h1;
            {4'h4, 5'h3}: color = 5'h1;
            {4'h4, 5'h4}: color = 5'h1;
            {4'h4, 5'h5}: color = 5'h2;
            {4'h4, 5'h6}: color = 5'h2;
            {4'h4, 5'h7}: color = 5'h2;
            {4'h4, 5'h8}: color = 5'h3;
            {4'h4, 5'h9}: color = 5'h3;
            {4'h4, 5'hA}: color = 5'h3;
            {4'h4, 5'hB}: color = 5'h3;
            {4'h4, 5'hC}: color = 5'h4;
            {4'h4, 5'hD}: color = 5'h4;
            {4'h4, 5'hE}: color = 5'h4;
            {4'h4, 5'hF}: color = 5'h5;
            {4'h4, 5'h10}: color = 5'h5;
            {4'h4, 5'h11}: color = 5'h5;
            {4'h4, 5'h12}: color = 5'h6;
            {4'h4, 5'h13}: color = 5'h6;
            {4'h4, 5'h14}: color = 5'h6;
            {4'h4, 5'h15}: color = 5'h7;
            {4'h4, 5'h16}: color = 5'h7;
            {4'h4, 5'h17}: color = 5'h7;
            {4'h4, 5'h18}: color = 5'h8;
            {4'h4, 5'h19}: color = 5'h8;
            {4'h4, 5'h1A}: color = 5'h8;
            {4'h4, 5'h1B}: color = 5'h8;
            {4'h4, 5'h1C}: color = 5'h9;
            {4'h4, 5'h1D}: color = 5'h9;
            {4'h4, 5'h1E}: color = 5'h9;
            {4'h4, 5'h1F}: color = 5'hA;
            {4'h5, 5'h0}: color = 5'h0;
            {4'h5, 5'h1}: color = 5'h0;
            {4'h5, 5'h2}: color = 5'h1;
            {4'h5, 5'h3}: color = 5'h1;
            {4'h5, 5'h4}: color = 5'h2;
            {4'h5, 5'h5}: color = 5'h2;
            {4'h5, 5'h6}: color = 5'h2;
            {4'h5, 5'h7}: color = 5'h3;
            {4'h5, 5'h8}: color = 5'h3;
            {4'h5, 5'h9}: color = 5'h3;
            {4'h5, 5'hA}: color = 5'h4;
            {4'h5, 5'hB}: color = 5'h4;
            {4'h5, 5'hC}: color = 5'h5;
            {4'h5, 5'hD}: color = 5'h5;
            {4'h5, 5'hE}: color = 5'h5;
            {4'h5, 5'hF}: color = 5'h6;
            {4'h5, 5'h10}: color = 5'h6;
            {4'h5, 5'h11}: color = 5'h6;
            {4'h5, 5'h12}: color = 5'h7;
            {4'h5, 5'h13}: color = 5'h7;
            {4'h5, 5'h14}: color = 5'h8;
            {4'h5, 5'h15}: color = 5'h8;
            {4'h5, 5'h16}: color = 5'h8;
            {4'h5, 5'h17}: color = 5'h9;
            {4'h5, 5'h18}: color = 5'h9;
            {4'h5, 5'h19}: color = 5'h9;
            {4'h5, 5'h1A}: color = 5'hA;
            {4'h5, 5'h1B}: color = 5'hA;
            {4'h5, 5'h1C}: color = 5'hB;
            {4'h5, 5'h1D}: color = 5'hB;
            {4'h5, 5'h1E}: color = 5'hB;
            {4'h5, 5'h1F}: color = 5'hC;
            {4'h6, 5'h0}: color = 5'h0;
            {4'h6, 5'h1}: color = 5'h0;
            {4'h6, 5'h2}: color = 5'h1;
            {4'h6, 5'h3}: color = 5'h1;
            {4'h6, 5'h4}: color = 5'h2;
            {4'h6, 5'h5}: color = 5'h2;
            {4'h6, 5'h6}: color = 5'h3;
            {4'h6, 5'h7}: color = 5'h3;
            {4'h6, 5'h8}: color = 5'h4;
            {4'h6, 5'h9}: color = 5'h4;
            {4'h6, 5'hA}: color = 5'h4;
            {4'h6, 5'hB}: color = 5'h5;
            {4'h6, 5'hC}: color = 5'h5;
            {4'h6, 5'hD}: color = 5'h6;
            {4'h6, 5'hE}: color = 5'h6;
            {4'h6, 5'hF}: color = 5'h7;
            {4'h6, 5'h10}: color = 5'h7;
            {4'h6, 5'h11}: color = 5'h7;
            {4'h6, 5'h12}: color = 5'h8;
            {4'h6, 5'h13}: color = 5'h8;
            {4'h6, 5'h14}: color = 5'h9;
            {4'h6, 5'h15}: color = 5'h9;
            {4'h6, 5'h16}: color = 5'hA;
            {4'h6, 5'h17}: color = 5'hA;
            {4'h6, 5'h18}: color = 5'hB;
            {4'h6, 5'h19}: color = 5'hB;
            {4'h6, 5'h1A}: color = 5'hB;
            {4'h6, 5'h1B}: color = 5'hC;
            {4'h6, 5'h1C}: color = 5'hC;
            {4'h6, 5'h1D}: color = 5'hD;
            {4'h6, 5'h1E}: color = 5'hD;
            {4'h6, 5'h1F}: color = 5'hE;
            {4'h7, 5'h0}: color = 5'h0;
            {4'h7, 5'h1}: color = 5'h1;
            {4'h7, 5'h2}: color = 5'h1;
            {4'h7, 5'h3}: color = 5'h2;
            {4'h7, 5'h4}: color = 5'h2;
            {4'h7, 5'h5}: color = 5'h3;
            {4'h7, 5'h6}: color = 5'h3;
            {4'h7, 5'h7}: color = 5'h4;
            {4'h7, 5'h8}: color = 5'h4;
            {4'h7, 5'h9}: color = 5'h5;
            {4'h7, 5'hA}: color = 5'h5;
            {4'h7, 5'hB}: color = 5'h6;
            {4'h7, 5'hC}: color = 5'h6;
            {4'h7, 5'hD}: color = 5'h7;
            {4'h7, 5'hE}: color = 5'h7;
            {4'h7, 5'hF}: color = 5'h8;
            {4'h7, 5'h10}: color = 5'h8;
            {4'h7, 5'h11}: color = 5'h9;
            {4'h7, 5'h12}: color = 5'h9;
            {4'h7, 5'h13}: color = 5'hA;
            {4'h7, 5'h14}: color = 5'hA;
            {4'h7, 5'h15}: color = 5'hB;
            {4'h7, 5'h16}: color = 5'hB;
            {4'h7, 5'h17}: color = 5'hC;
            {4'h7, 5'h18}: color = 5'hC;
            {4'h7, 5'h19}: color = 5'hD;
            {4'h7, 5'h1A}: color = 5'hD;
            {4'h7, 5'h1B}: color = 5'hE;
            {4'h7, 5'h1C}: color = 5'hE;
            {4'h7, 5'h1D}: color = 5'hF;
            {4'h7, 5'h1E}: color = 5'hF;
            {4'h7, 5'h1F}: color = 5'h10;
            {4'h8, 5'h0}: color = 5'h0;
            {4'h8, 5'h1}: color = 5'h1;
            {4'h8, 5'h2}: color = 5'h1;
            {4'h8, 5'h3}: color = 5'h2;
            {4'h8, 5'h4}: color = 5'h2;
            {4'h8, 5'h5}: color = 5'h3;
            {4'h8, 5'h6}: color = 5'h3;
            {4'h8, 5'h7}: color = 5'h4;
            {4'h8, 5'h8}: color = 5'h5;
            {4'h8, 5'h9}: color = 5'h5;
            {4'h8, 5'hA}: color = 5'h6;
            {4'h8, 5'hB}: color = 5'h6;
            {4'h8, 5'hC}: color = 5'h7;
            {4'h8, 5'hD}: color = 5'h7;
            {4'h8, 5'hE}: color = 5'h8;
            {4'h8, 5'hF}: color = 5'h8;
            {4'h8, 5'h10}: color = 5'h9;
            {4'h8, 5'h11}: color = 5'hA;
            {4'h8, 5'h12}: color = 5'hA;
            {4'h8, 5'h13}: color = 5'hB;
            {4'h8, 5'h14}: color = 5'hB;
            {4'h8, 5'h15}: color = 5'hC;
            {4'h8, 5'h16}: color = 5'hC;
            {4'h8, 5'h17}: color = 5'hD;
            {4'h8, 5'h18}: color = 5'hE;
            {4'h8, 5'h19}: color = 5'hE;
            {4'h8, 5'h1A}: color = 5'hF;
            {4'h8, 5'h1B}: color = 5'hF;
            {4'h8, 5'h1C}: color = 5'h10;
            {4'h8, 5'h1D}: color = 5'h10;
            {4'h8, 5'h1E}: color = 5'h11;
            {4'h8, 5'h1F}: color = 5'h11;
            {4'h9, 5'h0}: color = 5'h0;
            {4'h9, 5'h1}: color = 5'h1;
            {4'h9, 5'h2}: color = 5'h1;
            {4'h9, 5'h3}: color = 5'h2;
            {4'h9, 5'h4}: color = 5'h3;
            {4'h9, 5'h5}: color = 5'h3;
            {4'h9, 5'h6}: color = 5'h4;
            {4'h9, 5'h7}: color = 5'h4;
            {4'h9, 5'h8}: color = 5'h5;
            {4'h9, 5'h9}: color = 5'h6;
            {4'h9, 5'hA}: color = 5'h6;
            {4'h9, 5'hB}: color = 5'h7;
            {4'h9, 5'hC}: color = 5'h8;
            {4'h9, 5'hD}: color = 5'h8;
            {4'h9, 5'hE}: color = 5'h9;
            {4'h9, 5'hF}: color = 5'h9;
            {4'h9, 5'h10}: color = 5'hA;
            {4'h9, 5'h11}: color = 5'hB;
            {4'h9, 5'h12}: color = 5'hB;
            {4'h9, 5'h13}: color = 5'hC;
            {4'h9, 5'h14}: color = 5'hD;
            {4'h9, 5'h15}: color = 5'hD;
            {4'h9, 5'h16}: color = 5'hE;
            {4'h9, 5'h17}: color = 5'hE;
            {4'h9, 5'h18}: color = 5'hF;
            {4'h9, 5'h19}: color = 5'h10;
            {4'h9, 5'h1A}: color = 5'h10;
            {4'h9, 5'h1B}: color = 5'h11;
            {4'h9, 5'h1C}: color = 5'h12;
            {4'h9, 5'h1D}: color = 5'h12;
            {4'h9, 5'h1E}: color = 5'h13;
            {4'h9, 5'h1F}: color = 5'h13;
            {4'hA, 5'h0}: color = 5'h0;
            {4'hA, 5'h1}: color = 5'h1;
            {4'hA, 5'h2}: color = 5'h1;
            {4'hA, 5'h3}: color = 5'h2;
            {4'hA, 5'h4}: color = 5'h3;
            {4'hA, 5'h5}: color = 5'h3;
            {4'hA, 5'h6}: color = 5'h4;
            {4'hA, 5'h7}: color = 5'h5;
            {4'hA, 5'h8}: color = 5'h6;
            {4'hA, 5'h9}: color = 5'h6;
            {4'hA, 5'hA}: color = 5'h7;
            {4'hA, 5'hB}: color = 5'h8;
            {4'hA, 5'hC}: color = 5'h8;
            {4'hA, 5'hD}: color = 5'h9;
            {4'hA, 5'hE}: color = 5'hA;
            {4'hA, 5'hF}: color = 5'hA;
            {4'hA, 5'h10}: color = 5'hB;
            {4'hA, 5'h11}: color = 5'hC;
            {4'hA, 5'h12}: color = 5'hC;
            {4'hA, 5'h13}: color = 5'hD;
            {4'hA, 5'h14}: color = 5'hE;
            {4'hA, 5'h15}: color = 5'hE;
            {4'hA, 5'h16}: color = 5'hF;
            {4'hA, 5'h17}: color = 5'h10;
            {4'hA, 5'h18}: color = 5'h11;
            {4'hA, 5'h19}: color = 5'h11;
            {4'hA, 5'h1A}: color = 5'h12;
            {4'hA, 5'h1B}: color = 5'h13;
            {4'hA, 5'h1C}: color = 5'h13;
            {4'hA, 5'h1D}: color = 5'h14;
            {4'hA, 5'h1E}: color = 5'h15;
            {4'hA, 5'h1F}: color = 5'h15;
            {4'hB, 5'h0}: color = 5'h0;
            {4'hB, 5'h1}: color = 5'h1;
            {4'hB, 5'h2}: color = 5'h2;
            {4'hB, 5'h3}: color = 5'h2;
            {4'hB, 5'h4}: color = 5'h3;
            {4'hB, 5'h5}: color = 5'h4;
            {4'hB, 5'h6}: color = 5'h5;
            {4'hB, 5'h7}: color = 5'h5;
            {4'hB, 5'h8}: color = 5'h6;
            {4'hB, 5'h9}: color = 5'h7;
            {4'hB, 5'hA}: color = 5'h8;
            {4'hB, 5'hB}: color = 5'h8;
            {4'hB, 5'hC}: color = 5'h9;
            {4'hB, 5'hD}: color = 5'hA;
            {4'hB, 5'hE}: color = 5'hB;
            {4'hB, 5'hF}: color = 5'hB;
            {4'hB, 5'h10}: color = 5'hC;
            {4'hB, 5'h11}: color = 5'hD;
            {4'hB, 5'h12}: color = 5'hE;
            {4'hB, 5'h13}: color = 5'hE;
            {4'hB, 5'h14}: color = 5'hF;
            {4'hB, 5'h15}: color = 5'h10;
            {4'hB, 5'h16}: color = 5'h11;
            {4'hB, 5'h17}: color = 5'h11;
            {4'hB, 5'h18}: color = 5'h12;
            {4'hB, 5'h19}: color = 5'h13;
            {4'hB, 5'h1A}: color = 5'h14;
            {4'hB, 5'h1B}: color = 5'h14;
            {4'hB, 5'h1C}: color = 5'h15;
            {4'hB, 5'h1D}: color = 5'h16;
            {4'hB, 5'h1E}: color = 5'h17;
            {4'hB, 5'h1F}: color = 5'h17;
            {4'hC, 5'h0}: color = 5'h0;
            {4'hC, 5'h1}: color = 5'h1;
            {4'hC, 5'h2}: color = 5'h2;
            {4'hC, 5'h3}: color = 5'h2;
            {4'hC, 5'h4}: color = 5'h3;
            {4'hC, 5'h5}: color = 5'h4;
            {4'hC, 5'h6}: color = 5'h5;
            {4'hC, 5'h7}: color = 5'h6;
            {4'hC, 5'h8}: color = 5'h7;
            {4'hC, 5'h9}: color = 5'h7;
            {4'hC, 5'hA}: color = 5'h8;
            {4'hC, 5'hB}: color = 5'h9;
            {4'hC, 5'hC}: color = 5'hA;
            {4'hC, 5'hD}: color = 5'hB;
            {4'hC, 5'hE}: color = 5'hB;
            {4'hC, 5'hF}: color = 5'hC;
            {4'hC, 5'h10}: color = 5'hD;
            {4'hC, 5'h11}: color = 5'hE;
            {4'hC, 5'h12}: color = 5'hF;
            {4'hC, 5'h13}: color = 5'hF;
            {4'hC, 5'h14}: color = 5'h10;
            {4'hC, 5'h15}: color = 5'h11;
            {4'hC, 5'h16}: color = 5'h12;
            {4'hC, 5'h17}: color = 5'h13;
            {4'hC, 5'h18}: color = 5'h14;
            {4'hC, 5'h19}: color = 5'h14;
            {4'hC, 5'h1A}: color = 5'h15;
            {4'hC, 5'h1B}: color = 5'h16;
            {4'hC, 5'h1C}: color = 5'h17;
            {4'hC, 5'h1D}: color = 5'h18;
            {4'hC, 5'h1E}: color = 5'h18;
            {4'hC, 5'h1F}: color = 5'h19;
            {4'hD, 5'h0}: color = 5'h0;
            {4'hD, 5'h1}: color = 5'h1;
            {4'hD, 5'h2}: color = 5'h2;
            {4'hD, 5'h3}: color = 5'h3;
            {4'hD, 5'h4}: color = 5'h4;
            {4'hD, 5'h5}: color = 5'h4;
            {4'hD, 5'h6}: color = 5'h5;
            {4'hD, 5'h7}: color = 5'h6;
            {4'hD, 5'h8}: color = 5'h7;
            {4'hD, 5'h9}: color = 5'h8;
            {4'hD, 5'hA}: color = 5'h9;
            {4'hD, 5'hB}: color = 5'hA;
            {4'hD, 5'hC}: color = 5'hB;
            {4'hD, 5'hD}: color = 5'hB;
            {4'hD, 5'hE}: color = 5'hC;
            {4'hD, 5'hF}: color = 5'hD;
            {4'hD, 5'h10}: color = 5'hE;
            {4'hD, 5'h11}: color = 5'hF;
            {4'hD, 5'h12}: color = 5'h10;
            {4'hD, 5'h13}: color = 5'h11;
            {4'hD, 5'h14}: color = 5'h12;
            {4'hD, 5'h15}: color = 5'h12;
            {4'hD, 5'h16}: color = 5'h13;
            {4'hD, 5'h17}: color = 5'h14;
            {4'hD, 5'h18}: color = 5'h15;
            {4'hD, 5'h19}: color = 5'h16;
            {4'hD, 5'h1A}: color = 5'h17;
            {4'hD, 5'h1B}: color = 5'h18;
            {4'hD, 5'h1C}: color = 5'h19;
            {4'hD, 5'h1D}: color = 5'h19;
            {4'hD, 5'h1E}: color = 5'h1A;
            {4'hD, 5'h1F}: color = 5'h1B;
            {4'hE, 5'h0}: color = 5'h0;
            {4'hE, 5'h1}: color = 5'h1;
            {4'hE, 5'h2}: color = 5'h2;
            {4'hE, 5'h3}: color = 5'h3;
            {4'hE, 5'h4}: color = 5'h4;
            {4'hE, 5'h5}: color = 5'h5;
            {4'hE, 5'h6}: color = 5'h6;
            {4'hE, 5'h7}: color = 5'h7;
            {4'hE, 5'h8}: color = 5'h8;
            {4'hE, 5'h9}: color = 5'h8;
            {4'hE, 5'hA}: color = 5'h9;
            {4'hE, 5'hB}: color = 5'hA;
            {4'hE, 5'hC}: color = 5'hB;
            {4'hE, 5'hD}: color = 5'hC;
            {4'hE, 5'hE}: color = 5'hD;
            {4'hE, 5'hF}: color = 5'hE;
            {4'hE, 5'h10}: color = 5'hF;
            {4'hE, 5'h11}: color = 5'h10;
            {4'hE, 5'h12}: color = 5'h11;
            {4'hE, 5'h13}: color = 5'h12;
            {4'hE, 5'h14}: color = 5'h13;
            {4'hE, 5'h15}: color = 5'h14;
            {4'hE, 5'h16}: color = 5'h15;
            {4'hE, 5'h17}: color = 5'h16;
            {4'hE, 5'h18}: color = 5'h17;
            {4'hE, 5'h19}: color = 5'h17;
            {4'hE, 5'h1A}: color = 5'h18;
            {4'hE, 5'h1B}: color = 5'h19;
            {4'hE, 5'h1C}: color = 5'h1A;
            {4'hE, 5'h1D}: color = 5'h1B;
            {4'hE, 5'h1E}: color = 5'h1C;
            {4'hE, 5'h1F}: color = 5'h1D;
            {4'hF, 5'h0}: color = 5'h0;
            {4'hF, 5'h1}: color = 5'h1;
            {4'hF, 5'h2}: color = 5'h2;
            {4'hF, 5'h3}: color = 5'h3;
            {4'hF, 5'h4}: color = 5'h4;
            {4'hF, 5'h5}: color = 5'h5;
            {4'hF, 5'h6}: color = 5'h6;
            {4'hF, 5'h7}: color = 5'h7;
            {4'hF, 5'h8}: color = 5'h8;
            {4'hF, 5'h9}: color = 5'h9;
            {4'hF, 5'hA}: color = 5'hA;
            {4'hF, 5'hB}: color = 5'hB;
            {4'hF, 5'hC}: color = 5'hC;
            {4'hF, 5'hD}: color = 5'hD;
            {4'hF, 5'hE}: color = 5'hE;
            {4'hF, 5'hF}: color = 5'hF;
            {4'hF, 5'h10}: color = 5'h10;
            {4'hF, 5'h11}: color = 5'h11;
            {4'hF, 5'h12}: color = 5'h12;
            {4'hF, 5'h13}: color = 5'h13;
            {4'hF, 5'h14}: color = 5'h14;
            {4'hF, 5'h15}: color = 5'h15;
            {4'hF, 5'h16}: color = 5'h16;
            {4'hF, 5'h17}: color = 5'h17;
            {4'hF, 5'h18}: color = 5'h18;
            {4'hF, 5'h19}: color = 5'h19;
            {4'hF, 5'h1A}: color = 5'h1A;
            {4'hF, 5'h1B}: color = 5'h1B;
            {4'hF, 5'h1C}: color = 5'h1C;
            {4'hF, 5'h1D}: color = 5'h1D;
            {4'hF, 5'h1E}: color = 5'h1E;
            {4'hF, 5'h1F}: color = 5'h1F;
            default: color = 5'h0;
        endcase
    end
    
endmodule
